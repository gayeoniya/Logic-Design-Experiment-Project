// [���� �߰���] ��ư ��ٿ�� ��� (Array ����)
module Debounce_Array #(
    parameter WIDTH = 8
)(
    input wire clk,
    input wire rst_n,
    input wire [WIDTH-1:0] btn_in,
    output reg [WIDTH-1:0] btn_out
);

    // 50MHz Ŭ�� ����, �� 20ms ��ٿ��
    // 20ms / 20ns = 1,000,000 count
    localparam CNT_MAX = 1000000;

    reg [WIDTH-1:0] btn_prev;
    reg [19:0] cnt [WIDTH-1:0]; // �� ��ư�� ī����
    
    genvar i;
    generate
        for (i = 0; i < WIDTH; i = i + 1) begin : db_loop
            always @(posedge clk or negedge rst_n) begin
                if (!rst_n) begin
                    cnt[i] <= 0;
                    btn_out[i] <= 0;
                    btn_prev[i] <= 0;
                end else begin
                    // �Է� ���°� �������� ī���� ����
                    if (btn_in[i] != btn_prev[i]) begin
                        cnt[i] <= 0;
                        btn_prev[i] <= btn_in[i];
                    end else if (cnt[i] < CNT_MAX) begin
                        cnt[i] <= cnt[i] + 1;
                    end else begin
                        // ���� �ð� �����Ǹ� ��� ������Ʈ
                        btn_out[i] <= btn_prev[i];
                    end
                end
            end
        end
    endgenerate

endmodule

// ���� ��Ʈ�� (Start ��ư��)
module Debounce (
    input wire clk,
    input wire rst_n,
    input wire btn_in,
    output reg btn_out
);
    localparam CNT_MAX = 1000000; // 20ms
    reg btn_prev;
    reg [19:0] cnt;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            cnt <= 0;
            btn_out <= 0;
            btn_prev <= 0;
        end else begin
            if (btn_in != btn_prev) begin
                cnt <= 0;
                btn_prev <= btn_in;
            end else if (cnt < CNT_MAX) begin
                cnt <= cnt + 1;
            end else begin
                btn_out <= btn_prev;
            end
        end
    end
endmodule
module LCD_Display_Controller (
    input wire clk,             // 50MHz Clock
    input wire rst_n,
    input wire [127:0] line_1,  // LCD ù° �� ������ (16����)
    input wire [127:0] line_2,  // LCD ��° �� ������ (16����)

    // ���� LCD�� ������ ��ȣ (Top ����� Output�� ��)
    output reg lcd_rs,          // 0: ���, 1: ������
    output reg lcd_rw,          // 0: ���� (�׻� 0)
    output reg lcd_en,          // Enable ��ȣ
    output reg [7:0] lcd_data   // 8��Ʈ ������ ����
);

    // ���� ����
    localparam S_IDLE       = 4'd0;
    localparam S_INIT       = 4'd1;  // �ʱ�ȭ
    localparam S_LINE1      = 4'd2;  // ù° �� ��� ��
    localparam S_LINE2      = 4'd3;  // ��° �� ��� ��
    localparam S_DELAY      = 4'd4;  // ��� ó�� ���

    reg [3:0] state;
    reg [3:0] next_state;
    
    // [����] �ռ� ������ ���·� �ʱ�ȭ ��ɾ� ó��
    // initial ��� �����ϰ� case������ ó��
    
    reg [2:0] init_idx;      // �ʱ�ȭ �ܰ� ī����
    reg [3:0] char_idx;      // ���� ���� ī���� (0~15)
    reg [19:0] delay_cnt;    // ������ ī����
    
    // 50MHz ���� ������ ����
    localparam DELAY_TIME = 100000; 

    // �ʱ�ȭ ��ɾ� ���� �Լ� (Combinational)
    function [7:0] get_init_cmd;
        input [2:0] idx;
        begin
            case (idx)
                3'd0: get_init_cmd = 8'h38; // 8-bit mode, 2 lines
                3'd1: get_init_cmd = 8'h0C; // Display ON, Cursor OFF
                3'd2: get_init_cmd = 8'h06; // Auto Increment
                3'd3: get_init_cmd = 8'h01; // Clear Display
                3'd4: get_init_cmd = 8'h80; // Cursor Home
                default: get_init_cmd = 8'h00;
            endcase
        end
    endfunction

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= S_INIT;
            init_idx <= 0;
            char_idx <= 0;
            lcd_en <= 0;
            lcd_rs <= 0;
            lcd_rw <= 0;
            lcd_data <= 0;
            delay_cnt <= 0;
        end else begin
            case (state)
                // 1. �ʱ�ȭ �ܰ�
                S_INIT: begin
                    lcd_rs <= 0; // ��� ���
                    lcd_rw <= 0;
                    lcd_data <= get_init_cmd(init_idx); // �Լ� ȣ��� ����
                    
                    if (delay_cnt == 0) lcd_en <= 1; // Pulse High
                    if (delay_cnt == 5000) lcd_en <= 0; // Pulse Low (Enable �� Ȯ��)
                    
                    if (delay_cnt < DELAY_TIME) begin
                        delay_cnt <= delay_cnt + 1;
                    end else begin
                        delay_cnt <= 0;
                        if (init_idx < 4) begin
                            init_idx <= init_idx + 1;
                        end else begin
                            state <= S_LINE1; // �ʱ�ȭ ��, ��� ����
                            char_idx <= 0;
                        end
                    end
                end

                // 2. ù ��° �� ���
                S_LINE1: begin
                    lcd_rs <= 1; // ������ ��� (���� ����)
                    lcd_rw <= 0;
                    
                    // 128��Ʈ �����Ϳ��� �ش� ����(char_idx)�� ����(8��Ʈ) �̾Ƴ���
                    lcd_data <= line_1[127 - (char_idx * 8) -: 8];

                    if (delay_cnt == 0) lcd_en <= 1;
                    if (delay_cnt == 2000) lcd_en <= 0;

                    if (delay_cnt < 5000) begin 
                        delay_cnt <= delay_cnt + 1;
                    end else begin
                        delay_cnt <= 0;
                        if (char_idx < 15) begin
                            char_idx <= char_idx + 1;
                        end else begin
                            // �� �ٲ� �غ� (Ŀ���� �� ��° �ٷ� �̵�: 0xC0)
                            state <= S_DELAY;
                            next_state <= S_LINE2;
                            lcd_rs <= 0; // ���
                            lcd_data <= 8'hC0; 
                        end
                    end
                end

                // 3. �� �ٲ� �� �߰� ��� ó��
                S_DELAY: begin
                      if (delay_cnt == 0) lcd_en <= 1;
                      if (delay_cnt == 5000) lcd_en <= 0;
                      
                      if (delay_cnt < DELAY_TIME) delay_cnt <= delay_cnt + 1;
                      else begin
                          delay_cnt <= 0;
                          state <= next_state;
                          char_idx <= 0;
                      end
                end

                // 4. �� ��° �� ���
                S_LINE2: begin
                    lcd_rs <= 1; 
                    lcd_data <= line_2[127 - (char_idx * 8) -: 8];

                    if (delay_cnt == 0) lcd_en <= 1;
                    if (delay_cnt == 2000) lcd_en <= 0;

                    if (delay_cnt < 5000) begin
                        delay_cnt <= delay_cnt + 1;
                    end else begin
                        delay_cnt <= 0;
                        if (char_idx < 15) begin
                            char_idx <= char_idx + 1;
                        end else begin
                            // �ٽ� ó������ (Ŀ�� Ȩ: 0x80)
                            state <= S_DELAY;
                            next_state <= S_LINE1; // ��� ����
                            lcd_rs <= 0;
                            lcd_data <= 8'h80;
                        end
                    end
                end
            endcase
        end
    end
endmodule
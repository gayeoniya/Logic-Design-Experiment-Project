module Display_7Seg (
    input clk,
    input rst_n,
    input [31:0] user_seq,      
    input [3:0] input_cnt,      
    
    output reg [7:0] seg_data,
    output reg [7:0] seg_sel    
);
    reg [19:0] scan_cnt;
    wire [2:0] scan_idx;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) scan_cnt <= 20'd0;
        else        scan_cnt <= scan_cnt + 1;
    end
    
    // ��ĵ �ӵ� ����
    assign scan_idx = scan_cnt[19:17];

    reg [3:0] display_num;
    
    always @(*) begin
        // �⺻������ ��� �� (Active Low ���� 11111111)
        seg_sel = 8'hFF; 
        display_num = 4'd15; // 15 = Blank (Empty)

        // [������] Digit 0(���� ������ ��)���� 1, 2, 3... ������ ä�������� ����
        case (scan_idx)
            // 0��° �ڸ� (Digit 0) -> ù ��° �Է°� ǥ��
            3'd0: begin 
                seg_sel = ~8'b00000001; 
                if (input_cnt >= 1) display_num = user_seq[3:0];
            end
            
            // 1��° �ڸ� (Digit 1) -> �� ��° �Է°� ǥ��
            3'd1: begin 
                seg_sel = ~8'b00000010;
                if (input_cnt >= 2) display_num = user_seq[7:4];
            end
            
            // 2��° �ڸ� (Digit 2) -> �� ��° �Է°� ǥ��
            3'd2: begin 
                seg_sel = ~8'b00000100;
                if (input_cnt >= 3) display_num = user_seq[11:8];
            end
            
            // 3��° �ڸ� (Digit 3) -> �� ��° �Է°� ǥ��
            3'd3: begin 
                seg_sel = ~8'b00001000;
                if (input_cnt >= 4) display_num = user_seq[15:12];
            end
            
            // 4��° �ڸ� (Digit 4) -> �ټ� ��° �Է°� ǥ��
            3'd4: begin 
                seg_sel = ~8'b00010000;
                if (input_cnt >= 5) display_num = user_seq[19:16];
            end
            
            // 5��° �ڸ� (Digit 5) -> ���� ��° �Է°� ǥ��
            3'd5: begin 
                seg_sel = ~8'b00100000;
                if (input_cnt >= 6) display_num = user_seq[23:20];
            end
            
            // 6��° �ڸ� (Digit 6) -> �ϰ� ��° �Է°� ǥ��
            3'd6: begin 
                seg_sel = ~8'b01000000;
                if (input_cnt >= 7) display_num = user_seq[27:24];
            end
            
            // 7��° �ڸ� (Digit 7) -> ���� ��° �Է°� ǥ��
            3'd7: begin 
                seg_sel = ~8'b10000000;
                if (input_cnt >= 8) display_num = user_seq[31:28];
            end
        endcase
    end

    reg [7:0] decode_out;
    always @(*) begin
        case (display_num)
            // ���� ���� ���� (0�� ���� ����)
            4'd0: decode_out = 8'b1100_0000; 
            4'd1: decode_out = 8'b1111_1001;
            4'd2: decode_out = 8'b1010_0100;
            4'd3: decode_out = 8'b1011_0000;
            4'd4: decode_out = 8'b1001_1001;
            4'd5: decode_out = 8'b1001_0010;
            4'd6: decode_out = 8'b1000_0010;
            4'd7: decode_out = 8'b1111_1000;
            4'd8: decode_out = 8'b1000_0000;
            4'd9: decode_out = 8'b1001_0000;
            default: decode_out = 8'b1111_1111; // OFF
        endcase
        
        // [������] ȹ�� �ݴ�� ���´ٸ� ������ ��ȣ�� �������Ѿ� �մϴ�.
        // ���� �ڵ忡�� ~�� �߰��Ͽ� �������׽��ϴ�.
        seg_data = ~decode_out; 
    end
endmodule
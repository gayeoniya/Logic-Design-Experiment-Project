module LCD_Text_Gen (
    input [2:0] state,            // FSM ����
    input [2:0] current_round,    // ���� ����
    input [15:0] total_score,     // ���� ����
    input is_success,             // ���� ���� (S_PASS �� 1)

    // LCD�� ���� ������ (16���� * 8��Ʈ = 128��Ʈ)
    output reg [127:0] line_1,    
    output reg [127:0] line_2     
);

    // ====================================================
    // 1. ���ڸ� ASCII �ڵ�� ��ȯ (0~9 -> '0'~'9')
    // ====================================================
    wire [7:0] ascii_round;
    wire [7:0] ascii_score_100, ascii_score_10, ascii_score_1;

    // ���� ��ȯ
    assign ascii_round = {5'd0, current_round} + 8'h30;
    
    // ���� ��ȯ (100�� �ڸ�, 10�� �ڸ�, 1�� �ڸ�)
    assign ascii_score_100 = ((total_score / 100) % 10) + 8'h30;
    assign ascii_score_10  = ((total_score / 10) % 10)  + 8'h30;
    assign ascii_score_1   = (total_score % 10)         + 8'h30;

    // ====================================================
    // 2. FSM ���°� ���� (Game_FSM�� ����)
    // ====================================================
    localparam S_IDLE       = 3'd0;
    localparam S_GEN_SEQ    = 3'd1; 
    localparam S_SHOW_SEQ   = 3'd2; 
    localparam S_WAIT_INPUT = 3'd3;
    localparam S_CHECK      = 3'd4; 
    localparam S_PASS       = 3'd5;
    localparam S_FAIL       = 3'd6; 
    localparam S_DONE       = 3'd7;

    // ====================================================
    // 3. LCD ��� �ؽ�Ʈ ���� ����
    // ====================================================
    always @(*) begin
        // [�߿�] Latch ������ ���� �⺻ �ʱ�ȭ (��� ����)
        line_1 = "                "; 
        line_2 = "                ";

        case (state)
            // ---------------------------------------------------------
            // [ȭ�� 1] ���� ��� ȭ��
            // ---------------------------------------------------------
            S_IDLE: begin
                line_1 = "   Game Start   "; 
                line_2 = "                ";
            end

            // ---------------------------------------------------------
            // [ȭ�� 2] ���� �÷��� ȭ�� (���� / ���� ǥ��)
            // �� ������: S_CHECK ���¸� ���⿡ ���Խ��׽��ϴ�.
            // ���� Ȯ�� ��� �ð�(0.5��) ���� ���� ȭ���� �����Ͽ�
            // ����� ������ ���� "Fail..."�� �����̴� ������ �����ϴ�.
            // ---------------------------------------------------------
            S_GEN_SEQ, S_SHOW_SEQ, S_WAIT_INPUT, S_CHECK: begin
                // Line 1: "Lv. 1           "
                line_1[127:96] = "Lv. ";  
                line_1[95:88]  = ascii_round; 

                // Line 2: "Score: 000      "
                line_2[127:72] = "Score: "; 
                line_2[71:64]  = ascii_score_100;
                line_2[63:56]  = ascii_score_10; 
                line_2[55:48]  = ascii_score_1;  
            end

            // ---------------------------------------------------------
            // [ȭ�� 3] ���� ��� ȭ�� (����/����)
            // ���� ����� Ȯ���� S_PASS, S_FAIL������ ������ ���ϴ�.
            // ---------------------------------------------------------
            S_PASS, S_FAIL: begin
                if (state == S_FAIL) begin
                    // ���� ��
                    line_1 = "     Fail...    ";
                    line_2 = "  Try Again...  ";
                end else begin
                    // ���� �� (S_PASS)
                    line_1 = "    Success!    ";
                    line_2 = " Next Level...  ";
                end
            end

            // ---------------------------------------------------------
            // [ȭ�� 4] ���� ���� Ŭ���� (��� ���� ����)
            // ---------------------------------------------------------
            S_DONE: begin
                line_1 = "  FINAL SCORE   ";
                // Line 2: "  Total: 100    "
                line_2[127:72] = "    Total: ";
                line_2[71:64]  = ascii_score_100;
                line_2[63:56]  = ascii_score_10;
                line_2[55:48]  = ascii_score_1;
            end
            
            // ---------------------------------------------------------
            // ���� ó��
            // ---------------------------------------------------------
            default: begin
                line_1 = "   System Err   ";
                line_2 = "  Check State   ";
            end
        endcase
    end

endmodule